module alu_control(opcode,cadd, cflag_out,calu_out,op_adder,op_logic,op_bitops,add_size);
input [5:0]opcode;
output [2:0] cflag_out;
output [1:0] calu_out;
output op_adder;
output [1:0] op_logic;
output [2:0] op_bitops;
output [1:0] cadd;
output add_size;
reg [1:0] cadd;
reg [2:0] cflag_out;
reg [1:0] calu_out;
reg op_adder;
reg [1:0] op_logic;
reg [2:0] op_bitops;
reg add_size;

always@(opcode)
begin
	case(opcode)
	6'h00:begin//add
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b00;
				add_size=1'b0;
				op_logic=2'b0;
				op_bitops=3'b0;
				end
	6'h01:begin//addi
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b01;
				add_size=1'b0;
				op_logic=2'b0;
				op_bitops=3'b0;
				end
	6'h02:begin//sub
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b1;
				cadd=2'b00;
				add_size=1'b0;
				op_logic=2'b0;
				op_bitops=3'b0;
				end
	6'h03:begin//add16
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b00;
				add_size=1'b1;
				op_logic=2'b0;
				op_bitops=3'b0;
				end
	6'h04:begin//addi16
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b01;
				add_size=1'b1;
				op_logic=2'b0;
				op_bitops=3'b0;
				end
	6'h05:begin//sub16
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b1;
				cadd=2'b00;
				add_size=1'b1;
				op_logic=2'b0;
				op_bitops=3'b0;
				end
	6'h1a:begin//subi
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b1;
				cadd=2'b01;
				add_size=1'b0;
				op_logic=2'b0;
				op_bitops=3'b0;
				end
	6'h1b:begin//subi16
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b1;
				cadd=2'b01;
				add_size=1'b1;
				op_logic=2'b0;
				op_bitops=3'b0;
				end
	6'h06:begin//and
				cflag_out=3'b010;
				calu_out=2'b10;
				op_logic=2'b00;
				cadd=2'b00;
				op_adder=1'b0;
				op_bitops=3'b0;
				add_size=1'b0;
				end
	6'h07:begin//andi
				cflag_out=3'b010;
				op_adder=1'b0;
				op_logic=2'b00;
				cadd=2'b01;
				calu_out=2'b10;
				op_bitops=3'b0;
				add_size=1'b0;
				end
	6'h08:begin//or
				cflag_out=3'b010;
				calu_out=2'b10;
				op_logic=2'b01;
				cadd=2'b00;
				op_adder=1'b0;
				op_bitops=3'b0;
				add_size=1'b0;
				end
	6'h09:begin//ori
				cflag_out=3'b010;
				calu_out=2'b10;
				op_logic=2'b01;
				cadd=2'b01;
				op_adder=1'b0;
				op_bitops=3'b0;
				add_size=1'b0;
				end
	6'h0a:begin//xor
				cflag_out=3'b010;
				calu_out=2'b10;
				op_logic=2'b10;
				cadd=2'b00;
				op_adder=1'b0;
				op_bitops=3'b0;
				add_size=1'b0;
				end
	6'h0b:begin//xori
				cflag_out=3'b010;
				calu_out=2'b10;
				op_logic=2'b10;
				cadd=2'b01;
				op_adder=1'b0;
				op_bitops=3'b0;
				add_size=1'b0;
				end
	6'h0c:begin//not
				cflag_out=3'b010;
				calu_out=2'b10;
				op_logic=2'b11;
				cadd=2'b00;
				op_adder=1'b0;
				op_bitops=3'b0;
				add_size=1'b0;
				end
	6'h0d:begin//shiftrotate
				cflag_out=3'b011;
				calu_out=2'b11;
				op_logic=2'b00;
				op_adder=1'b0;
				op_bitops=3'b0;
				cadd=2'b0;
				add_size=1'b0;
				end
	6'h0e:begin//get4
				cflag_out=3'b001;
				calu_out=2'b01;
				op_bitops=3'b100;
				op_logic=2'b00;
				op_adder=1'b0;
				cadd=2'b0;
				add_size=1'b0;
				end
	6'h0f:begin//merge4
				cflag_out=3'b001;
				calu_out=2'b01;
				op_bitops=3'b101;
				op_logic=2'b00;
				op_adder=1'b0;
				cadd=2'b0;
				add_size=1'b0;
				end
	6'h11:begin//daa
				cflag_out=3'b100;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b10;
				add_size=1'b0;//adds in 8-bit may need 16 bit
				op_bitops=3'b000;
				op_logic=2'b00;
				end
	6'h12:begin//getbit
				cflag_out=3'b001;
				calu_out=2'b01;
				op_bitops=3'b000;
				op_logic=2'b00;
				op_adder=1'b0;
				cadd=2'b0;
				add_size=1'b0;
				end
	6'h13:begin//ngetbit
				cflag_out=3'b001;
				calu_out=2'b01;
				op_bitops=3'b001;
				op_logic=2'b00;
				op_adder=1'b0;
				cadd=2'b0;
				add_size=1'b0;
				end
	6'h14:begin//setbit
				cflag_out=3'b001;
				calu_out=2'b01;
				op_bitops=3'b010;
				op_logic=2'b00;
				op_adder=1'b0;
				cadd=2'b0;
				add_size=1'b0;
				end
	6'h15:begin//nsetbit
				cflag_out=3'b001;
				calu_out=2'b01;
				op_bitops=3'b011;
				op_logic=2'b00;
				op_adder=1'b0;
				cadd=2'b0;
				add_size=1'b0;
				end
	6'h30:begin//ld
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b01;
				add_size=1'b0;
				op_bitops=3'b000;
				op_logic=2'b00;
				end
	6'h31:begin//st
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b01;
				add_size=1'b0;
				op_bitops=3'b000;
				op_logic=2'b00;
				end
	6'h16:begin//limm
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b01;
				add_size=1'b1;
				op_bitops=3'b000;
				op_logic=2'b00;
				end
	6'h32:begin//in
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b01;
				add_size=1'b0;
				op_bitops=3'b000;
				op_logic=2'b00;
				end
	6'h33:begin//out
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				cadd=2'b01;
				add_size=1'b0;
				op_bitops=3'b000;
				op_logic=2'b00;
				end
	default:begin
				cflag_out=3'b000;
				calu_out=2'b00;
				op_adder=1'b0;
				op_logic=2'b00;
				op_bitops=3'b00;
				cadd=2'b00;
				add_size=1'b0;
				end
	endcase
end//always
endmodule